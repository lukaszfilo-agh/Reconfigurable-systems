`timescale 1ns / 1ps
//-----------------------------------------------
// Company: agh
//-----------------------------------------------
module i_mem
(
  input [7:0]address,
  output [31:0]data
);
//-----------------------------------------------
//instruction memory
wire [31:0]program[255:0];
//movi R1, 0x03
assign program[0] = 32'b00000000_00110000_10000001_00000011;
//movi R2, 0x60
assign program[1] = 32'b00000000_00110000_10000010_01100000;
//loadi R4, 0x6
assign program[2] = 32'b00000000_00110000_10001100_00000110;
//load R4, R1
assign program[3] = 32'b00000000_00010001_10001100_00000000;
//jz R4, 0x0C
assign program[4] = 32'b00000010_00110100_10000110_00001100;
//movi R5, 0xE1
assign program[5] = 32'b00000000_00110000_10000101_11100001;
//andi R5, R5, 0xD3
assign program[6] = 32'b00000000_00000101_10000101_11010011;
//add R3, R1, R2
assign program[7] = 32'b00000000_00010001_00100011_00000000;
//movi R2, 0x00
assign program[8] = 32'b00000000_00110000_10000010_00000000;
//add R0, R3, R1
assign program[9] = 32'b00000000_00010011_00010000_00000000;
//addi R1, R1, 0x01
assign program[10] = 32'b00000000_00010001_10000001_00000001;
//jumpi 0x02
assign program[11] = 32'b00000001_00110000_10000110_00000010;
//nop
assign program[12] = 32'b00000000_00000000_00000110_00000000;
//nop
assign program[13] = 32'b00000000_00000000_00000110_00000000;
//nop
assign program[14] = 32'b00000000_00000000_00000110_00000000;
//movi R1, 0x03
assign program[15] = 32'b00000000_00110000_10000001_00000011;
//jump R1
assign program[16] = 32'b00000001_00010001_10000110_00000000;


//// movi R0, 0x34
//assign program[0]= 32'b00000000_00010110_10000000_00110100;
//// mov R1, R0
//assign program[1]= 32'b00000000_00010000_01100001_00000000;
//// nop
//assign program[2]= 32'b00000000_00000000_00000110_00000000;


//-----------------------------------------------
assign data=program[address];
//-----------------------------------------------
endmodule
//-----------------------------------------------

`timescale 1ns / 1ps
//-----------------------------------------------
// Company: agh
//-----------------------------------------------
module i_mem
(
  input [7:0]address,
  output [31:0]data
);
//-----------------------------------------------
//instruction memory
wire [31:0]program[255:0];

//movi R4, 0x01
assign program[0] = 32'b00000000_00110000_10000100_00000001;
//movi R2, 0x22
assign program[1] = 32'b00000000_00110000_10000010_00100010;
//movi R1, 0x22
assign program[2] = 32'b00000000_00110000_10000001_00100010;
//movi R0, 0x22
assign program[3] = 32'b00000000_00110000_10000000_00100010;
//addi R0, R0, 0x01
assign program[4] = 32'b00000000_00010000_10000000_00000001;
//jnz R0, 0x04
assign program[5] = 32'b00000011_00110000_10000110_00000100;
//addi R1, R1, 0x01
assign program[6] = 32'b00000000_00010001_10000001_00000001;
//jnz R1, 0x04
assign program[7] = 32'b00000011_00110001_10000110_00000100;
//addi R2, R2, 0x01
assign program[8] = 32'b00000000_00010010_10000010_00000001;
//jnz R2, 0x04
assign program[9] = 32'b00000011_00110010_10000110_00000100;
//movi R2, 0x22
assign program[10] = 32'b00000000_00110000_10000010_00100010;
//movi R1, 0x22
assign program[11] = 32'b00000000_00110000_10000001_00100010;
//movi R0, 0x22
assign program[12] = 32'b00000000_00110000_10000000_00100010;
//addi R0, R0, 0x01
assign program[13] = 32'b00000000_00010000_10000000_00000001;
//jnz R0, 0x0D
assign program[14] = 32'b00000011_00110000_10000110_00001101;
//addi R1, R1, 0x01
assign program[15] = 32'b00000000_00010001_10000001_00000001;
//jnz R1, 0x0D
assign program[16] = 32'b00000011_00110001_10000110_00001101;
//addi R2, R2, 0x01
assign program[17] = 32'b00000000_00010010_10000010_00000001;
//jnz R2, 0x0D
assign program[18] = 32'b00000011_00110010_10000110_00001101;
//movi R4, 0x02
assign program[19] = 32'b00000000_00110000_10000100_00000010;
//andi R3, R5, 0x01
assign program[20] = 32'b00000000_00000101_10000011_00000001;
//jz R3, 0x14
assign program[21] = 32'b00000010_00110011_10000110_00010100;
//movi R4, 0x04
assign program[22] = 32'b00000000_00110000_10000100_00000100;
//movi R2, 0x22
assign program[23] = 32'b00000000_00110000_10000010_00100010;
//movi R1, 0x22
assign program[24] = 32'b00000000_00110000_10000001_00100010;
//movi R0, 0x22
assign program[25] = 32'b00000000_00110000_10000000_00100010;
//addi R0, R0, 0x01
assign program[26] = 32'b00000000_00010000_10000000_00000001;
//jnz R0, 0x1A
assign program[27] = 32'b00000011_00110000_10000110_00011010;
//addi R1, R1, 0x01
assign program[28] = 32'b00000000_00010001_10000001_00000001;
//jnz R1, 0x1A
assign program[29] = 32'b00000011_00110001_10000110_00011010;
//addi R2, R2, 0x01
assign program[30] = 32'b00000000_00010010_10000010_00000001;
//jnz R2, 0x1A
assign program[31] = 32'b00000011_00110010_10000110_00011010;
//movi R4, 0x04
assign program[32] = 32'b00000000_00110000_10000100_00000100;
//movi R2, 0x22
assign program[33] = 32'b00000000_00110000_10000010_00100010;
//movi R1, 0x22
assign program[34] = 32'b00000000_00110000_10000001_00100010;
//movi R0, 0x22
assign program[35] = 32'b00000000_00110000_10000000_00100010;
//addi R0, R0, 0x01
assign program[36] = 32'b00000000_00010000_10000000_00000001;
//jnz R0, 0x24
assign program[37] = 32'b00000011_00110000_10000110_00100100;
//addi R1, R1, 0x01
assign program[38] = 32'b00000000_00010001_10000001_00000001;
//jnz R1, 0x24
assign program[39] = 32'b00000011_00110001_10000110_00100100;
//addi R2, R2, 0x01
assign program[40] = 32'b00000000_00010010_10000010_00000001;
//jnz R2, 0x24
assign program[41] = 32'b00000011_00110010_10000110_00100100;
//movi R4, 0x08
assign program[42] = 32'b00000000_00110000_10000100_00001000;
//andi R3, R5, 0x02
assign program[43] = 32'b00000000_00000101_10000011_00000010;
//jz R3, 0x2B
assign program[44] = 32'b00000010_00110011_10000110_00101011;
//jumpi 0x00
assign program[45] = 32'b00000001_00110000_10000110_00000000;







//-----------------------------------------------
assign data=program[address];
//-----------------------------------------------
endmodule
//-----------------------------------------------
